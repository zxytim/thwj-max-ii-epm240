-- megafunction wizard: %ALTUFM_SPI%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTUFM_SPI 

-- ============================================================
-- File Name: altufm_spa.vhd
-- Megafunction Name(s):
-- 			ALTUFM_SPI
--
-- Simulation Library Files(s):
-- 			maxii
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 12.1 Build 243 01/31/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2012 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altufm_spi ACCESS_MODE="READ_ONLY" BYTE_OF_PAGE_WRITE=8 CBX_AUTO_BLACKBOX="ALL" CONFIG_MODE="BASE" DEVICE_FAMILY="MAX II" ERASE_TIME=500000000 LPM_FILE="data.hex" OSC_FREQUENCY=180000 PROGRAM_TIME=1600000 WIDTH_UFM_ADDRESS=9 ncs osc sck si so
--VERSION_BEGIN 12.1SP1 cbx_a_gray2bin 2013:01:31:18:04:54:SJ cbx_a_graycounter 2013:01:31:18:04:54:SJ cbx_altufm_spi 2013:01:31:18:04:55:SJ cbx_cycloneii 2013:01:31:18:04:55:SJ cbx_lpm_add_sub 2013:01:31:18:04:55:SJ cbx_lpm_compare 2013:01:31:18:04:55:SJ cbx_lpm_counter 2013:01:31:18:04:55:SJ cbx_lpm_decode 2013:01:31:18:04:55:SJ cbx_lpm_mux 2013:01:31:18:04:55:SJ cbx_maxii 2013:01:31:18:04:55:SJ cbx_mgl 2013:01:31:18:08:38:SJ cbx_stratix 2013:01:31:18:04:55:SJ cbx_stratixii 2013:01:31:18:04:55:SJ cbx_util_mgl 2013:01:31:18:04:55:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

 LIBRARY maxii;
 USE maxii.all;

--synthesis_resources = a_graycounter 3 lpm_counter 1 lut 55 maxii_ufm 1 TRI 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altufm_spa_altufm_spi_5bl IS 
	 PORT 
	 ( 
		 ncs	:	IN  STD_LOGIC;
		 osc	:	OUT  STD_LOGIC;
		 sck	:	IN  STD_LOGIC;
		 si	:	IN  STD_LOGIC;
		 so	:	OUT  STD_LOGIC
	 ); 
 END altufm_spa_altufm_spi_5bl;

 ARCHITECTURE RTL OF altufm_spa_altufm_spi_5bl IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c101;suppress_da_rule_internal=c103;suppress_da_rule_internal=c104;suppress_da_rule_internal=c106;suppress_da_rule_internal=d101;suppress_da_rule_internal=r101;suppress_da_rule_internal=s102;suppress_da_rule_internal=s104";

	 SIGNAL  wire_address_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_ncs_wire1w80w81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_cntr_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_data_cntr_w_lg_w_q_range93w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_data_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_ncs_wire1w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_data_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_data_cntr_w_q_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_cntr_w_lg_w_q_range10w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_cntr_w_lg_w_q_range8w9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_ncs_wire1w5w6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_op_cntr_w_q_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_cntr_w_q_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 addr_cmplt_dly	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 addr_cmplt_dly2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 addr_sload_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_addr_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_addr_dly_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_addr_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_addr_reg_ena	:	STD_LOGIC;
	 SIGNAL	 op_cmplt_dly	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 op_cnt_stage	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 op_cnt_stage2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 op_code7_dly	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_op_code7_dly_ena	:	STD_LOGIC;
	 SIGNAL  wire_op_code7_dly_w_lg_q186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_op_code_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 op_code_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_op_code_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_lg_w_lg_w_lg_w72w73w74w75w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_lg_w_lg_w72w73w74w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_lg_w72w73w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w72w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_lg_w_lg_w_lg_w_q_range67w68w69w70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_lg_w_lg_w_q_range67w68w69w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_lg_w_q_range67w68w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_q_range24w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_q_range27w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_q_range30w64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_q_range33w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_q_range36w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_lg_w_q_range67w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_op_code_reg_w_q_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_op_code_streg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 op_code_streg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_op_code_streg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_rd_addr_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 rd_addr_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_rd_addr_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_addr_sload133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_read_addr_cntr_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_maxii_ufm_block1_bgpbusy	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_busy	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_drdout	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_osc	:	STD_LOGIC;
	 SIGNAL	 wire_tri_buf2_out	:	STD_LOGIC;
	 SIGNAL	 wire_tri_buf2_oe	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_sck_wire182w183w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_ncs_wire1w15w16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sck_wire182w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_ncs_wire1w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_ncs_wire1w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_ncs_wire1w5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_op_complete104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sck_wire182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_complete_dly103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_address_complete79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data_complete190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_addr179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ncs_wire1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_op_complete2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_addr_lim127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sck_wire4w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ufm_bgpbusy14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ufm_busy61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  addr_complete_dly :	STD_LOGIC;
	 SIGNAL  addr_complete_dly2 :	STD_LOGIC;
	 SIGNAL  addr_sload :	STD_LOGIC;
	 SIGNAL  addr_to_cmplt :	STD_LOGIC;
	 SIGNAL  address_complete :	STD_LOGIC;
	 SIGNAL  circuit_reset :	STD_LOGIC;
	 SIGNAL  data_complete :	STD_LOGIC;
	 SIGNAL  end_addr :	STD_LOGIC;
	 SIGNAL  init_end_addr :	STD_LOGIC;
	 SIGNAL  ncs_wire :	STD_LOGIC;
	 SIGNAL  op_code7 :	STD_LOGIC;
	 SIGNAL  op_complete :	STD_LOGIC;
	 SIGNAL  op_complete_dly :	STD_LOGIC;
	 SIGNAL  op_stage :	STD_LOGIC;
	 SIGNAL  oscena	:	STD_LOGIC;
	 SIGNAL  reach_addr_lim :	STD_LOGIC;
	 SIGNAL  read_op :	STD_LOGIC;
	 SIGNAL  sck_wire :	STD_LOGIC;
	 SIGNAL  si_wire :	STD_LOGIC;
	 SIGNAL  so_wire :	STD_LOGIC;
	 SIGNAL  ufm_arclk :	STD_LOGIC;
	 SIGNAL  ufm_ardin :	STD_LOGIC;
	 SIGNAL  ufm_arshft :	STD_LOGIC;
	 SIGNAL  ufm_bgpbusy :	STD_LOGIC;
	 SIGNAL  ufm_busy :	STD_LOGIC;
	 SIGNAL  ufm_drclk :	STD_LOGIC;
	 SIGNAL  ufm_drdin :	STD_LOGIC;
	 SIGNAL  ufm_drdout :	STD_LOGIC;
	 SIGNAL  ufm_drshft :	STD_LOGIC;
	 SIGNAL  ufm_erase :	STD_LOGIC;
	 SIGNAL  ufm_osc :	STD_LOGIC;
	 SIGNAL  ufm_oscena :	STD_LOGIC;
	 SIGNAL  ufm_program :	STD_LOGIC;
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  maxii_ufm
	 GENERIC 
	 (
		ADDRESS_WIDTH	:	NATURAL := 9;
		ERASE_TIME	:	NATURAL := 500000000;
		INIT_FILE	:	STRING := "UNUSED";
		mem1	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem10	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem11	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem12	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem13	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem14	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem15	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem16	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem2	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem3	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem4	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem5	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem6	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem7	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem8	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem9	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		OSC_SIM_SETTING	:	NATURAL := 180000;
		PROGRAM_TIME	:	NATURAL := 1600000;
		lpm_type	:	STRING := "maxii_ufm"
	 );
	 PORT
	 ( 
		arclk	:	IN STD_LOGIC := '0';
		ardin	:	IN STD_LOGIC := '0';
		arshft	:	IN STD_LOGIC := '1';
		bgpbusy	:	OUT STD_LOGIC;
		busy	:	OUT STD_LOGIC;
		drclk	:	IN STD_LOGIC := '0';
		drdin	:	IN STD_LOGIC := '0';
		drdout	:	OUT STD_LOGIC;
		drshft	:	IN STD_LOGIC := '1';
		erase	:	IN STD_LOGIC := '0';
		osc	:	OUT STD_LOGIC;
		oscena	:	IN STD_LOGIC := '0';
		program	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_sck_wire182w183w184w(0) <= wire_w_lg_w_lg_sck_wire182w183w(0) AND read_op;
	wire_w_lg_w_lg_w_lg_ncs_wire1w15w16w(0) <= wire_w_lg_w_lg_ncs_wire1w15w(0) AND wire_w_lg_ufm_bgpbusy14w(0);
	wire_w_lg_w_lg_sck_wire182w183w(0) <= wire_w_lg_sck_wire182w(0) AND wire_w_lg_addr_complete_dly103w(0);
	wire_w_lg_w_lg_ncs_wire1w15w(0) <= wire_w_lg_ncs_wire1w(0) AND wire_w_lg_op_complete2w(0);
	wire_w_lg_w_lg_ncs_wire1w80w(0) <= wire_w_lg_ncs_wire1w(0) AND op_complete;
	wire_w_lg_w_lg_ncs_wire1w5w(0) <= wire_w_lg_ncs_wire1w(0) AND op_stage;
	wire_w_lg_op_complete104w(0) <= op_complete AND wire_w_lg_addr_complete_dly103w(0);
	wire_w_lg_sck_wire182w(0) <= sck_wire AND op_complete;
	wire_w_lg_addr_complete_dly103w(0) <= NOT addr_complete_dly;
	wire_w_lg_address_complete79w(0) <= NOT address_complete;
	wire_w_lg_data_complete190w(0) <= NOT data_complete;
	wire_w_lg_end_addr179w(0) <= NOT end_addr;
	wire_w_lg_ncs_wire1w(0) <= NOT ncs_wire;
	wire_w_lg_op_complete2w(0) <= NOT op_complete;
	wire_w_lg_reach_addr_lim127w(0) <= NOT reach_addr_lim;
	wire_w_lg_sck_wire4w(0) <= NOT sck_wire;
	wire_w_lg_ufm_bgpbusy14w(0) <= NOT ufm_bgpbusy;
	wire_w_lg_ufm_busy61w(0) <= NOT ufm_busy;
	addr_complete_dly <= addr_cmplt_dly;
	addr_complete_dly2 <= addr_cmplt_dly2;
	addr_sload <= addr_sload_reg;
	addr_to_cmplt <= ((((NOT wire_address_cntr_q(0)) AND (NOT wire_address_cntr_q(1))) AND wire_address_cntr_q(2)) AND (NOT wire_address_cntr_q(3)));
	address_complete <= ((((NOT wire_address_cntr_q(0)) AND (NOT wire_address_cntr_q(1))) AND wire_address_cntr_q(2)) AND wire_address_cntr_q(3));
	circuit_reset <= ncs_wire;
	data_complete <= (((NOT wire_data_cntr_q(0)) AND (NOT wire_data_cntr_q(1))) AND wire_data_cntr_q(2));
	end_addr <= end_addr_reg;
	init_end_addr <= (((((((rd_addr_reg(7) AND rd_addr_reg(6)) AND rd_addr_reg(5)) AND rd_addr_reg(4)) AND rd_addr_reg(3)) AND rd_addr_reg(2)) AND rd_addr_reg(1)) AND rd_addr_reg(0));
	ncs_wire <= ncs;
	op_code7 <= (wire_op_cntr_w_lg_w_q_range10w100w(0) AND wire_op_cntr_q(2));
	op_complete <= (((NOT wire_op_cntr_q(0)) AND wire_op_cntr_w_lg_w_q_range8w9w(0)) AND wire_op_cntr_q(2));
	op_complete_dly <= op_cmplt_dly;
	op_stage <= op_cnt_stage2;
	osc <= ufm_osc;
	oscena <= '1';
	reach_addr_lim <= (((((((wire_read_addr_cntr_q(7) AND wire_read_addr_cntr_q(6)) AND wire_read_addr_cntr_q(5)) AND wire_read_addr_cntr_q(4)) AND wire_read_addr_cntr_q(3)) AND wire_read_addr_cntr_q(2)) AND wire_read_addr_cntr_q(1)) AND wire_read_addr_cntr_q(0));
	read_op <= ((wire_op_code_reg_w_lg_w_lg_w_lg_w_lg_w72w73w74w75w76w(0) AND wire_w_lg_ufm_busy61w(0)) AND wire_w_lg_ufm_bgpbusy14w(0));
	sck_wire <= sck;
	si_wire <= si;
	so <= so_wire;
	so_wire <= wire_tri_buf2_out;
	ufm_arclk <= (wire_w_lg_w_lg_w_lg_sck_wire182w183w184w(0) OR (wire_data_cntr_w_lg_w_q_range93w180w(0) AND wire_w_lg_end_addr179w(0)));
	ufm_ardin <= (((si_wire AND op_complete_dly) AND wire_w_lg_addr_complete_dly103w(0)) AND wire_w_lg_ufm_bgpbusy14w(0));
	ufm_arshft <= (wire_op_code7_dly_w_lg_q186w(0) AND wire_w_lg_ufm_bgpbusy14w(0));
	ufm_bgpbusy <= wire_maxii_ufm_block1_bgpbusy;
	ufm_busy <= wire_maxii_ufm_block1_busy;
	ufm_drclk <= ((wire_w_lg_sck_wire4w(0) AND read_op) AND addr_complete_dly);
	ufm_drdin <= '0';
	ufm_drdout <= wire_maxii_ufm_block1_drdout;
	ufm_drshft <= ((addr_complete_dly2 AND wire_w_lg_data_complete190w(0)) AND read_op);
	ufm_erase <= '0';
	ufm_osc <= wire_maxii_ufm_block1_osc;
	ufm_oscena <= oscena;
	ufm_program <= '0';
	wire_address_cntr_clk_en <= wire_w_lg_w_lg_w_lg_ncs_wire1w80w81w(0);
	wire_w_lg_w_lg_w_lg_ncs_wire1w80w81w(0) <= wire_w_lg_w_lg_ncs_wire1w80w(0) AND wire_w_lg_address_complete79w(0);
	address_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 4
	  )
	  PORT MAP ( 
		aclr => circuit_reset,
		clk_en => wire_address_cntr_clk_en,
		clock => sck_wire,
		q => wire_address_cntr_q
	  );
	wire_data_cntr_w_lg_w_q_range93w180w(0) <= wire_data_cntr_w_q_range93w(0) AND read_op;
	wire_data_cntr_clk_en <= wire_w_lg_w_lg_ncs_wire1w175w(0);
	wire_w_lg_w_lg_ncs_wire1w175w(0) <= wire_w_lg_ncs_wire1w(0) AND addr_complete_dly2;
	wire_data_cntr_w_q_range93w(0) <= wire_data_cntr_q(2);
	data_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => circuit_reset,
		clk_en => wire_data_cntr_clk_en,
		clock => sck_wire,
		q => wire_data_cntr_q
	  );
	wire_op_cntr_w_lg_w_q_range10w100w(0) <= wire_op_cntr_w_q_range10w(0) AND wire_op_cntr_w_lg_w_q_range8w9w(0);
	wire_op_cntr_w_lg_w_q_range8w9w(0) <= NOT wire_op_cntr_w_q_range8w(0);
	wire_op_cntr_clk_en <= wire_w_lg_w_lg_w_lg_ncs_wire1w5w6w(0);
	wire_w_lg_w_lg_w_lg_ncs_wire1w5w6w(0) <= wire_w_lg_w_lg_ncs_wire1w5w(0) AND wire_w_lg_op_complete2w(0);
	wire_op_cntr_w_q_range10w(0) <= wire_op_cntr_q(0);
	wire_op_cntr_w_q_range8w(0) <= wire_op_cntr_q(1);
	op_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => circuit_reset,
		clk_en => wire_op_cntr_clk_en,
		clock => sck_wire,
		q => wire_op_cntr_q
	  );
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN addr_cmplt_dly <= '0';
		ELSIF (sck_wire = '0' AND sck_wire'event) THEN 
			IF (ncs_wire = '0') THEN addr_cmplt_dly <= address_complete;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN addr_cmplt_dly2 <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (ncs_wire = '0') THEN addr_cmplt_dly2 <= address_complete;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN addr_sload_reg <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (read_op = '1') THEN addr_sload_reg <= addr_to_cmplt;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN end_addr_dly_reg <= '0';
		ELSIF (sck_wire = '0' AND sck_wire'event) THEN 
			IF (wire_end_addr_dly_reg_ena = '1') THEN end_addr_dly_reg <= reach_addr_lim;
			END IF;
		END IF;
	END PROCESS;
	wire_end_addr_dly_reg_ena <= (read_op AND data_complete);
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN end_addr_reg <= '0';
		ELSIF (sck_wire = '0' AND sck_wire'event) THEN 
			IF (wire_end_addr_reg_ena = '1') THEN end_addr_reg <= (init_end_addr OR end_addr_dly_reg);
			END IF;
		END IF;
	END PROCESS;
	wire_end_addr_reg_ena <= (read_op AND data_complete);
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_cmplt_dly <= '0';
		ELSIF (sck_wire = '0' AND sck_wire'event) THEN 
			IF (ncs_wire = '0') THEN op_cmplt_dly <= op_complete;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_cnt_stage <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (ncs_wire = '0') THEN op_cnt_stage <= wire_w_lg_op_complete2w(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_cnt_stage2 <= '0';
		ELSIF (sck_wire = '0' AND sck_wire'event) THEN 
			IF (ncs_wire = '0') THEN op_cnt_stage2 <= op_cnt_stage;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code7_dly <= '0';
		ELSIF (sck_wire = '0' AND sck_wire'event) THEN 
			IF (wire_op_code7_dly_ena = '1') THEN op_code7_dly <= op_code7;
			END IF;
		END IF;
	END PROCESS;
	wire_op_code7_dly_ena <= (wire_w_lg_ncs_wire1w(0) AND op_code7);
	wire_op_code7_dly_w_lg_q186w(0) <= op_code7_dly AND wire_w_lg_addr_complete_dly103w(0);
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(0) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(0) = '1') THEN op_code_reg(0) <= wire_op_code_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(1) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(1) = '1') THEN op_code_reg(1) <= wire_op_code_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(2) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(2) = '1') THEN op_code_reg(2) <= wire_op_code_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(3) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(3) = '1') THEN op_code_reg(3) <= wire_op_code_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(4) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(4) = '1') THEN op_code_reg(4) <= wire_op_code_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(5) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(5) = '1') THEN op_code_reg(5) <= wire_op_code_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(6) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(6) = '1') THEN op_code_reg(6) <= wire_op_code_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_reg(7) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_reg_ena(7) = '1') THEN op_code_reg(7) <= wire_op_code_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_op_code_reg_d <= ( op_code_reg(6 DOWNTO 0) & si_wire);
	loop0 : FOR i IN 0 TO 7 GENERATE
		wire_op_code_reg_ena(i) <= wire_w_lg_w_lg_w_lg_ncs_wire1w15w16w(0);
	END GENERATE loop0;
	wire_op_code_reg_w_lg_w_lg_w_lg_w_lg_w72w73w74w75w76w(0) <= wire_op_code_reg_w_lg_w_lg_w_lg_w72w73w74w75w(0) AND op_complete;
	wire_op_code_reg_w_lg_w_lg_w_lg_w72w73w74w75w(0) <= wire_op_code_reg_w_lg_w_lg_w72w73w74w(0) AND wire_op_code_reg_w_q_range19w(0);
	wire_op_code_reg_w_lg_w_lg_w72w73w74w(0) <= wire_op_code_reg_w_lg_w72w73w(0) AND wire_op_code_reg_w_q_range21w(0);
	wire_op_code_reg_w_lg_w72w73w(0) <= wire_op_code_reg_w72w(0) AND wire_op_code_reg_w_lg_w_q_range24w62w(0);
	wire_op_code_reg_w72w(0) <= wire_op_code_reg_w_lg_w_lg_w_lg_w_lg_w_q_range67w68w69w70w71w(0) AND wire_op_code_reg_w_lg_w_q_range27w63w(0);
	wire_op_code_reg_w_lg_w_lg_w_lg_w_lg_w_q_range67w68w69w70w71w(0) <= wire_op_code_reg_w_lg_w_lg_w_lg_w_q_range67w68w69w70w(0) AND wire_op_code_reg_w_lg_w_q_range30w64w(0);
	wire_op_code_reg_w_lg_w_lg_w_lg_w_q_range67w68w69w70w(0) <= wire_op_code_reg_w_lg_w_lg_w_q_range67w68w69w(0) AND wire_op_code_reg_w_lg_w_q_range33w65w(0);
	wire_op_code_reg_w_lg_w_lg_w_q_range67w68w69w(0) <= wire_op_code_reg_w_lg_w_q_range67w68w(0) AND wire_op_code_reg_w_lg_w_q_range36w66w(0);
	wire_op_code_reg_w_lg_w_q_range24w62w(0) <= NOT wire_op_code_reg_w_q_range24w(0);
	wire_op_code_reg_w_lg_w_q_range27w63w(0) <= NOT wire_op_code_reg_w_q_range27w(0);
	wire_op_code_reg_w_lg_w_q_range30w64w(0) <= NOT wire_op_code_reg_w_q_range30w(0);
	wire_op_code_reg_w_lg_w_q_range33w65w(0) <= NOT wire_op_code_reg_w_q_range33w(0);
	wire_op_code_reg_w_lg_w_q_range36w66w(0) <= NOT wire_op_code_reg_w_q_range36w(0);
	wire_op_code_reg_w_lg_w_q_range67w68w(0) <= NOT wire_op_code_reg_w_q_range67w(0);
	wire_op_code_reg_w_q_range19w(0) <= op_code_reg(0);
	wire_op_code_reg_w_q_range21w(0) <= op_code_reg(1);
	wire_op_code_reg_w_q_range24w(0) <= op_code_reg(2);
	wire_op_code_reg_w_q_range27w(0) <= op_code_reg(3);
	wire_op_code_reg_w_q_range30w(0) <= op_code_reg(4);
	wire_op_code_reg_w_q_range33w(0) <= op_code_reg(5);
	wire_op_code_reg_w_q_range36w(0) <= op_code_reg(6);
	wire_op_code_reg_w_q_range67w(0) <= op_code_reg(7);
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(0) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(0) = '1') THEN op_code_streg(0) <= wire_op_code_streg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(1) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(1) = '1') THEN op_code_streg(1) <= wire_op_code_streg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(2) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(2) = '1') THEN op_code_streg(2) <= wire_op_code_streg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(3) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(3) = '1') THEN op_code_streg(3) <= wire_op_code_streg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(4) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(4) = '1') THEN op_code_streg(4) <= wire_op_code_streg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(5) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(5) = '1') THEN op_code_streg(5) <= wire_op_code_streg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(6) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(6) = '1') THEN op_code_streg(6) <= wire_op_code_streg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN op_code_streg(7) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_op_code_streg_ena(7) = '1') THEN op_code_streg(7) <= wire_op_code_streg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_op_code_streg_d <= ( op_code_streg(6 DOWNTO 0) & si_wire);
	loop1 : FOR i IN 0 TO 7 GENERATE
		wire_op_code_streg_ena(i) <= wire_w_lg_w_lg_ncs_wire1w15w(0);
	END GENERATE loop1;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(0) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(0) = '1') THEN rd_addr_reg(0) <= wire_rd_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(1) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(1) = '1') THEN rd_addr_reg(1) <= wire_rd_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(2) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(2) = '1') THEN rd_addr_reg(2) <= wire_rd_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(3) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(3) = '1') THEN rd_addr_reg(3) <= wire_rd_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(4) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(4) = '1') THEN rd_addr_reg(4) <= wire_rd_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(5) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(5) = '1') THEN rd_addr_reg(5) <= wire_rd_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(6) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(6) = '1') THEN rd_addr_reg(6) <= wire_rd_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (sck_wire, circuit_reset)
	BEGIN
		IF (circuit_reset = '1') THEN rd_addr_reg(7) <= '0';
		ELSIF (sck_wire = '1' AND sck_wire'event) THEN 
			IF (wire_rd_addr_reg_ena(7) = '1') THEN rd_addr_reg(7) <= wire_rd_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_rd_addr_reg_d <= ( rd_addr_reg(6 DOWNTO 0) & si_wire);
	loop2 : FOR i IN 0 TO 7 GENERATE
		wire_rd_addr_reg_ena(i) <= wire_w_lg_op_complete104w(0);
	END GENERATE loop2;
	wire_read_addr_cntr_clk_en <= wire_w_lg_addr_sload133w(0);
	wire_w_lg_addr_sload133w(0) <= addr_sload OR (((((read_op AND address_complete) AND wire_w_lg_reach_addr_lim127w(0)) AND wire_data_cntr_q(2)) AND wire_data_cntr_q(1)) AND (NOT wire_data_cntr_q(0)));
	wire_read_addr_cntr_clock <= wire_w_lg_sck_wire4w(0);
	wire_read_addr_cntr_data <= ( rd_addr_reg(7 DOWNTO 0));
	read_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 8
	  )
	  PORT MAP ( 
		aclr => circuit_reset,
		clk_en => wire_read_addr_cntr_clk_en,
		clock => wire_read_addr_cntr_clock,
		data => wire_read_addr_cntr_data,
		q => wire_read_addr_cntr_q,
		sload => addr_sload
	  );
	maxii_ufm_block1 :  maxii_ufm
	  GENERIC MAP (
		ADDRESS_WIDTH => 9,
		ERASE_TIME => 500000000,
		INIT_FILE => "data.hex",
		mem1 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000111111111000000011111111100000001111111110000000111111111101010101111111110101010111111111010101011111111101010101111111110101010111111111010101011111111101010101111111110101010111111110000000111111111000000011111111100000001111111110000000111111111",
		mem10 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem11 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem12 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem13 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem14 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem15 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem16 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem2 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem3 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem4 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem5 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem6 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem7 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem8 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		mem9 => "00000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111",
		OSC_SIM_SETTING => 180000,
		PROGRAM_TIME => 1600000
	  )
	  PORT MAP ( 
		arclk => ufm_arclk,
		ardin => ufm_ardin,
		arshft => ufm_arshft,
		bgpbusy => wire_maxii_ufm_block1_bgpbusy,
		busy => wire_maxii_ufm_block1_busy,
		drclk => ufm_drclk,
		drdin => ufm_drdin,
		drdout => wire_maxii_ufm_block1_drdout,
		drshft => ufm_drshft,
		erase => ufm_erase,
		osc => wire_maxii_ufm_block1_osc,
		oscena => ufm_oscena,
		program => ufm_program
	  );
	wire_tri_buf2_out <= ufm_drdout WHEN wire_tri_buf2_oe = '1' ELSE 'Z';
	wire_tri_buf2_oe <= (((read_op AND addr_complete_dly) AND wire_w_lg_end_addr179w(0)) AND wire_w_lg_ncs_wire1w(0));

 END RTL; --altufm_spa_altufm_spi_5bl
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altufm_spa IS
	PORT
	(
		ncs		: IN STD_LOGIC ;
		sck		: IN STD_LOGIC ;
		si		: IN STD_LOGIC ;
		osc		: OUT STD_LOGIC ;
		so		: OUT STD_LOGIC 
	);
END altufm_spa;


ARCHITECTURE RTL OF altufm_spa IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTUFM_SPI";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "access_mode=READ_ONLY;byte_of_page_write=8;config_mode=BASE;erase_time=500000000;intended_device_family=MAX II;lpm_file=data.hex;lpm_hint=UNUSED;lpm_type=altufm_spi;osc_frequency=180000;program_time=1600000;width_ufm_address=9;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;



	COMPONENT altufm_spa_altufm_spi_5bl
	PORT (
			ncs	: IN STD_LOGIC ;
			si	: IN STD_LOGIC ;
			so	: OUT STD_LOGIC ;
			osc	: OUT STD_LOGIC ;
			sck	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	so    <= sub_wire0;
	osc    <= sub_wire1;

	altufm_spa_altufm_spi_5bl_component : altufm_spa_altufm_spi_5bl
	PORT MAP (
		ncs => ncs,
		si => si,
		sck => sck,
		so => sub_wire0,
		osc => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX II"
-- Retrieval info: PRIVATE: OSC_PORT STRING "ON"
-- Retrieval info: CONSTANT: ACCESS_MODE STRING "READ_ONLY"
-- Retrieval info: CONSTANT: BYTE_OF_PAGE_WRITE NUMERIC "8"
-- Retrieval info: CONSTANT: CONFIG_MODE STRING "BASE"
-- Retrieval info: CONSTANT: ERASE_TIME NUMERIC "500000000"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX II"
-- Retrieval info: CONSTANT: LPM_FILE STRING "data.hex"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altufm_spi"
-- Retrieval info: CONSTANT: OSC_FREQUENCY NUMERIC "180000"
-- Retrieval info: CONSTANT: PROGRAM_TIME NUMERIC "1600000"
-- Retrieval info: CONSTANT: WIDTH_UFM_ADDRESS NUMERIC "9"
-- Retrieval info: USED_PORT: ncs 0 0 0 0 INPUT NODEFVAL "ncs"
-- Retrieval info: CONNECT: @ncs 0 0 0 0 ncs 0 0 0 0
-- Retrieval info: USED_PORT: osc 0 0 0 0 OUTPUT NODEFVAL "osc"
-- Retrieval info: CONNECT: osc 0 0 0 0 @osc 0 0 0 0
-- Retrieval info: USED_PORT: sck 0 0 0 0 INPUT NODEFVAL "sck"
-- Retrieval info: CONNECT: @sck 0 0 0 0 sck 0 0 0 0
-- Retrieval info: USED_PORT: si 0 0 0 0 INPUT NODEFVAL "si"
-- Retrieval info: CONNECT: @si 0 0 0 0 si 0 0 0 0
-- Retrieval info: USED_PORT: so 0 0 0 0 OUTPUT NODEFVAL "so"
-- Retrieval info: CONNECT: so 0 0 0 0 @so 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altufm_spi.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altufm_spi.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altufm_spi.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altufm_spi_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altufm_spi.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altufm_spi.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: maxii
