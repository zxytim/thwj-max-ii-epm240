mem_spi_inst : mem_spi PORT MAP (
		ncs	 => ncs_sig,
		sck	 => sck_sig,
		si	 => si_sig,
		osc	 => osc_sig,
		so	 => so_sig
	);
