-- megafunction wizard: %ALTUFM_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTUFM_PARALLEL 

-- ============================================================
-- File Name: para.vhd
-- Megafunction Name(s):
-- 			ALTUFM_PARALLEL
--
-- Simulation Library Files(s):
-- 			maxii
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 12.1 Build 243 01/31/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2012 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altufm_parallel ACCESS_MODE="READ_ONLY" CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="MAX II" ERASE_TIME=500000000 OSC_FREQUENCY=180000 PROGRAM_TIME=1600000 WIDTH_ADDRESS=9 WIDTH_DATA=16 WIDTH_UFM_ADDRESS=9 addr data_valid dataout nbusy nread osc
--VERSION_BEGIN 12.1SP1 cbx_a_gray2bin 2013:01:31:18:04:54:SJ cbx_a_graycounter 2013:01:31:18:04:54:SJ cbx_altufm_parallel 2013:01:31:18:04:55:SJ cbx_cycloneii 2013:01:31:18:04:55:SJ cbx_lpm_add_sub 2013:01:31:18:04:55:SJ cbx_lpm_compare 2013:01:31:18:04:55:SJ cbx_lpm_counter 2013:01:31:18:04:55:SJ cbx_lpm_decode 2013:01:31:18:04:55:SJ cbx_lpm_mux 2013:01:31:18:04:55:SJ cbx_maxii 2013:01:31:18:04:55:SJ cbx_mgl 2013:01:31:18:08:38:SJ cbx_stratix 2013:01:31:18:04:55:SJ cbx_stratixii 2013:01:31:18:04:55:SJ cbx_util_mgl 2013:01:31:18:04:55:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

 LIBRARY maxii;
 USE maxii.all;

--synthesis_resources = lpm_counter 1 lut 62 maxii_ufm 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  para_altufm_parallel_t9l IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 data_valid	:	OUT  STD_LOGIC;
		 dataout	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 nbusy	:	OUT  STD_LOGIC;
		 nread	:	IN  STD_LOGIC;
		 osc	:	OUT  STD_LOGIC
	 ); 
 END para_altufm_parallel_t9l;

 ARCHITECTURE RTL OF para_altufm_parallel_t9l IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c101;suppress_da_rule_internal=c103;suppress_da_rule_internal=c104;suppress_da_rule_internal=r101;suppress_da_rule_internal=s104;suppress_da_rule_internal=s102";

	 SIGNAL	 A	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 data_valid_out_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 data_valid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_data_valid_reg_w_lg_q53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 deco1_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 decode_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 gated_clk1_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 gated_clk2_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 real_decode2_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_real_decode2_dffe_w_lg_q14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 real_decode_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sipo_dffe	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_tmp_do_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 tmp_do	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_tmp_do_ena	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
	 SIGNAL  wire_cntr2_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_maxii_ufm_block1_bgpbusy	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_drdout	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_osc	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_control_mux9w10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q224w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q335w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q335w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q335w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q44w25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr76w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_control_mux8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shiftin75w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_load74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_control_mux9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data_valid_en7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dly_tmp_decode17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nread1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tmp_decode52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ufm_bgpbusy12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ufm_osc165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q335w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_q335w36w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_q32w3w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_q32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_en :	STD_LOGIC;
	 SIGNAL  add_load :	STD_LOGIC;
	 SIGNAL  arclk :	STD_LOGIC;
	 SIGNAL  busy_arclk :	STD_LOGIC;
	 SIGNAL  busy_drclk :	STD_LOGIC;
	 SIGNAL  control_mux :	STD_LOGIC;
	 SIGNAL  copy_tmp_decode :	STD_LOGIC;
	 SIGNAL  data_valid_en :	STD_LOGIC;
	 SIGNAL  dly_tmp_decode :	STD_LOGIC;
	 SIGNAL  drdin :	STD_LOGIC;
	 SIGNAL  gated1 :	STD_LOGIC;
	 SIGNAL  gated2 :	STD_LOGIC;
	 SIGNAL  hold_decode :	STD_LOGIC;
	 SIGNAL  in_read_data_en :	STD_LOGIC;
	 SIGNAL  in_read_drclk :	STD_LOGIC;
	 SIGNAL  in_read_drshft :	STD_LOGIC;
	 SIGNAL  mux_nread :	STD_LOGIC;
	 SIGNAL  oscena	:	STD_LOGIC;
	 SIGNAL  q0 :	STD_LOGIC;
	 SIGNAL  q1 :	STD_LOGIC;
	 SIGNAL  q2 :	STD_LOGIC;
	 SIGNAL  q3 :	STD_LOGIC;
	 SIGNAL  q4 :	STD_LOGIC;
	 SIGNAL  read :	STD_LOGIC;
	 SIGNAL  read_op :	STD_LOGIC;
	 SIGNAL  real_decode :	STD_LOGIC;
	 SIGNAL  shiftin :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  sipo_q :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  start_decode :	STD_LOGIC;
	 SIGNAL  start_op :	STD_LOGIC;
	 SIGNAL  stop_op :	STD_LOGIC;
	 SIGNAL  tmp_add_en :	STD_LOGIC;
	 SIGNAL  tmp_add_load :	STD_LOGIC;
	 SIGNAL  tmp_arclk :	STD_LOGIC;
	 SIGNAL  tmp_arclk0 :	STD_LOGIC;
	 SIGNAL  tmp_ardin :	STD_LOGIC;
	 SIGNAL  tmp_arshft :	STD_LOGIC;
	 SIGNAL  tmp_data_valid2 :	STD_LOGIC;
	 SIGNAL  tmp_decode :	STD_LOGIC;
	 SIGNAL  tmp_drclk :	STD_LOGIC;
	 SIGNAL  tmp_in_read_data_en :	STD_LOGIC;
	 SIGNAL  tmp_in_read_drclk :	STD_LOGIC;
	 SIGNAL  tmp_in_read_drshft :	STD_LOGIC;
	 SIGNAL  tmp_read :	STD_LOGIC;
	 SIGNAL  ufm_arclk :	STD_LOGIC;
	 SIGNAL  ufm_ardin :	STD_LOGIC;
	 SIGNAL  ufm_arshft :	STD_LOGIC;
	 SIGNAL  ufm_bgpbusy :	STD_LOGIC;
	 SIGNAL  ufm_drclk :	STD_LOGIC;
	 SIGNAL  ufm_drdin :	STD_LOGIC;
	 SIGNAL  ufm_drdout :	STD_LOGIC;
	 SIGNAL  ufm_drshft :	STD_LOGIC;
	 SIGNAL  ufm_osc :	STD_LOGIC;
	 SIGNAL  ufm_oscena :	STD_LOGIC;
	 SIGNAL  X_var :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  Y_var :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  Z_var :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  maxii_ufm
	 GENERIC 
	 (
		ADDRESS_WIDTH	:	NATURAL := 9;
		ERASE_TIME	:	NATURAL := 500000000;
		INIT_FILE	:	STRING := "UNUSED";
		mem1	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem10	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem11	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem12	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem13	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem14	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem15	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem16	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem2	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem3	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem4	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem5	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem6	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem7	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem8	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem9	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		OSC_SIM_SETTING	:	NATURAL := 180000;
		PROGRAM_TIME	:	NATURAL := 1600000;
		lpm_type	:	STRING := "maxii_ufm"
	 );
	 PORT
	 ( 
		arclk	:	IN STD_LOGIC := '0';
		ardin	:	IN STD_LOGIC := '0';
		arshft	:	IN STD_LOGIC := '1';
		bgpbusy	:	OUT STD_LOGIC;
		busy	:	OUT STD_LOGIC;
		drclk	:	IN STD_LOGIC := '0';
		drdin	:	IN STD_LOGIC := '0';
		drdout	:	OUT STD_LOGIC;
		drshft	:	IN STD_LOGIC := '1';
		erase	:	IN STD_LOGIC := '0';
		osc	:	OUT STD_LOGIC;
		oscena	:	IN STD_LOGIC := '0';
		program	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_control_mux9w10w(0) <= wire_w_lg_control_mux9w(0) AND read;
	wire_w_lg_w_lg_q224w34w(0) <= wire_w_lg_q224w(0) AND wire_w_lg_q133w(0);
	wire_w_lg_w_lg_q335w59w(0) <= wire_w_lg_q335w(0) AND q0;
	wire_w_lg_w_lg_q335w58w(0) <= wire_w_lg_q335w(0) AND q1;
	wire_w_lg_w_lg_q335w60w(0) <= wire_w_lg_q335w(0) AND q2;
	wire_w_lg_w_lg_q44w25w(0) <= wire_w_lg_q44w(0) AND q3;
	loop0 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_addr76w(i) <= addr(i) AND add_load;
	END GENERATE loop0;
	wire_w_lg_control_mux8w(0) <= control_mux AND wire_w_lg_data_valid_en7w(0);
	wire_w_lg_q132w(0) <= q1 AND wire_w_lg_q031w(0);
	wire_w_lg_q356w(0) <= q3 AND wire_w_lg_q224w(0);
	wire_w_lg_q438w(0) <= q4 AND wire_w_lg_w_lg_w_lg_q335w36w37w(0);
	loop1 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_shiftin75w(i) <= shiftin(i) AND wire_w_lg_add_load74w(0);
	END GENERATE loop1;
	wire_w_lg_add_load74w(0) <= NOT add_load;
	wire_w_lg_control_mux9w(0) <= NOT control_mux;
	wire_w_lg_data_valid_en7w(0) <= NOT data_valid_en;
	wire_w_lg_dly_tmp_decode17w(0) <= NOT dly_tmp_decode;
	wire_w_lg_nread1w(0) <= NOT nread;
	wire_w_lg_q031w(0) <= NOT q0;
	wire_w_lg_q133w(0) <= NOT q1;
	wire_w_lg_q224w(0) <= NOT q2;
	wire_w_lg_q335w(0) <= NOT q3;
	wire_w_lg_q44w(0) <= NOT q4;
	wire_w_lg_tmp_decode52w(0) <= NOT tmp_decode;
	wire_w_lg_ufm_bgpbusy12w(0) <= NOT ufm_bgpbusy;
	wire_w_lg_ufm_osc165w(0) <= NOT ufm_osc;
	wire_w_lg_w_lg_q335w36w(0) <= wire_w_lg_q335w(0) OR wire_w_lg_w_lg_q224w34w(0);
	wire_w_lg_w_lg_w_lg_q335w36w37w(0) <= wire_w_lg_w_lg_q335w36w(0) OR wire_w_lg_q132w(0);
	wire_w_lg_w_lg_q32w3w(0) <= wire_w_lg_q32w(0) OR q1;
	wire_w_lg_q32w(0) <= q3 OR q2;
	add_en <= (tmp_add_en AND read_op);
	add_load <= (tmp_add_load AND read_op);
	arclk <= (tmp_arclk0 AND read_op);
	busy_arclk <= arclk;
	busy_drclk <= in_read_drclk;
	control_mux <= ((wire_w_lg_q44w(0) AND wire_w_lg_w_lg_q32w3w(0)) OR q4);
	copy_tmp_decode <= tmp_decode;
	data_valid <= data_valid_out_reg;
	data_valid_en <= ((q4 AND q3) AND q1);
	dataout <= tmp_do;
	dly_tmp_decode <= decode_dffe;
	drdin <= '0';
	gated1 <= gated_clk1_dffe;
	gated2 <= gated_clk2_dffe;
	hold_decode <= (wire_real_decode2_dffe_w_lg_q14w(0) AND real_decode);
	in_read_data_en <= (tmp_in_read_data_en AND read_op);
	in_read_drclk <= (tmp_in_read_drclk AND read_op);
	in_read_drshft <= (tmp_in_read_drshft AND read_op);
	mux_nread <= (wire_w_lg_w_lg_control_mux9w10w(0) OR wire_w_lg_control_mux8w(0));
	nbusy <= (wire_w_lg_dly_tmp_decode17w(0) AND wire_w_lg_ufm_bgpbusy12w(0));
	osc <= ufm_osc;
	oscena <= '1';
	q0 <= wire_cntr2_q(0);
	q1 <= wire_cntr2_q(1);
	q2 <= wire_cntr2_q(2);
	q3 <= wire_cntr2_q(3);
	q4 <= wire_cntr2_q(4);
	read <= wire_w_lg_nread1w(0);
	read_op <= tmp_read;
	real_decode <= start_decode;
	shiftin <= ( A(7 DOWNTO 0) & "0");
	sipo_q <= ( sipo_dffe(15 DOWNTO 0));
	start_decode <= (mux_nread AND wire_w_lg_ufm_bgpbusy12w(0));
	start_op <= (hold_decode OR stop_op);
	stop_op <= ((((q4 AND q3) AND wire_w_lg_q224w(0)) AND q1) AND q0);
	tmp_add_en <= (wire_w_lg_q44w(0) AND wire_w_lg_w_lg_q335w36w(0));
	tmp_add_load <= (NOT (wire_w_lg_q44w(0) AND (((wire_w_lg_w_lg_q335w60w(0) OR wire_w_lg_w_lg_q335w59w(0)) OR wire_w_lg_w_lg_q335w58w(0)) OR (wire_w_lg_q356w(0) AND wire_w_lg_q133w(0)))));
	tmp_arclk <= (gated1 AND wire_w_lg_ufm_osc165w(0));
	tmp_arclk0 <= (wire_w_lg_q44w(0) AND (wire_w_lg_q335w(0) OR (wire_w_lg_w_lg_q224w34w(0) AND wire_w_lg_q031w(0))));
	tmp_ardin <= A(8);
	tmp_arshft <= add_en;
	tmp_data_valid2 <= (stop_op AND read_op);
	tmp_decode <= tmp_read;
	tmp_drclk <= (gated2 AND wire_w_lg_ufm_osc165w(0));
	tmp_in_read_data_en <= ((wire_w_lg_q44w(0) AND ((q3 AND q2) OR (q3 AND q1))) OR wire_w_lg_q438w(0));
	tmp_in_read_drclk <= ((wire_w_lg_q44w(0) AND ((q3 AND q2) OR (q3 AND q1))) OR wire_w_lg_q438w(0));
	tmp_in_read_drshft <= (NOT (((wire_w_lg_w_lg_q44w25w(0) AND wire_w_lg_q224w(0)) AND q1) AND q0));
	tmp_read <= deco1_dffe;
	ufm_arclk <= tmp_arclk;
	ufm_ardin <= tmp_ardin;
	ufm_arshft <= tmp_arshft;
	ufm_bgpbusy <= wire_maxii_ufm_block1_bgpbusy;
	ufm_drclk <= tmp_drclk;
	ufm_drdin <= drdin;
	ufm_drdout <= wire_maxii_ufm_block1_drdout;
	ufm_drshft <= in_read_drshft;
	ufm_osc <= wire_maxii_ufm_block1_osc;
	ufm_oscena <= oscena;
	X_var <= wire_w_lg_shiftin75w;
	Y_var <= wire_w_lg_addr76w;
	Z_var <= (X_var OR Y_var);
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (add_en = '1') THEN A <= ( Z_var);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN data_valid_out_reg <= wire_data_valid_reg_w_lg_q53w(0);
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (data_valid_en = '1') THEN data_valid_reg <= tmp_data_valid2;
			END IF;
		END IF;
	END PROCESS;
	wire_data_valid_reg_w_lg_q53w(0) <= data_valid_reg AND wire_w_lg_tmp_decode52w(0);
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (start_op = '1') THEN deco1_dffe <= mux_nread;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN decode_dffe <= copy_tmp_decode;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN gated_clk1_dffe <= busy_arclk;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN gated_clk2_dffe <= busy_drclk;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN real_decode2_dffe <= real_decode_dffe;
		END IF;
	END PROCESS;
	wire_real_decode2_dffe_w_lg_q14w(0) <= NOT real_decode2_dffe;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN real_decode_dffe <= start_decode;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (in_read_data_en = '1') THEN sipo_dffe <= ( sipo_q(14 DOWNTO 0) & ufm_drdout);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(0) = '1') THEN tmp_do(0) <= wire_tmp_do_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(1) = '1') THEN tmp_do(1) <= wire_tmp_do_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(2) = '1') THEN tmp_do(2) <= wire_tmp_do_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(3) = '1') THEN tmp_do(3) <= wire_tmp_do_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(4) = '1') THEN tmp_do(4) <= wire_tmp_do_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(5) = '1') THEN tmp_do(5) <= wire_tmp_do_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(6) = '1') THEN tmp_do(6) <= wire_tmp_do_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(7) = '1') THEN tmp_do(7) <= wire_tmp_do_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(8) = '1') THEN tmp_do(8) <= wire_tmp_do_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(9) = '1') THEN tmp_do(9) <= wire_tmp_do_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(10) = '1') THEN tmp_do(10) <= wire_tmp_do_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(11) = '1') THEN tmp_do(11) <= wire_tmp_do_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(12) = '1') THEN tmp_do(12) <= wire_tmp_do_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(13) = '1') THEN tmp_do(13) <= wire_tmp_do_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(14) = '1') THEN tmp_do(14) <= wire_tmp_do_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (ufm_osc)
	BEGIN
		IF (ufm_osc = '1' AND ufm_osc'event) THEN 
			IF (wire_tmp_do_ena(15) = '1') THEN tmp_do(15) <= wire_tmp_do_d(15);
			END IF;
		END IF;
	END PROCESS;
	wire_tmp_do_d <= ( sipo_q(15 DOWNTO 0));
	loop2 : FOR i IN 0 TO 15 GENERATE
		wire_tmp_do_ena(i) <= wire_data_valid_reg_w_lg_q53w(0);
	END GENERATE loop2;
	cntr2 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_modulus => 28,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clk_en => tmp_decode,
		clock => ufm_osc,
		q => wire_cntr2_q
	  );
	maxii_ufm_block1 :  maxii_ufm
	  GENERIC MAP (
		ADDRESS_WIDTH => 9,
		ERASE_TIME => 500000000,
		INIT_FILE => "none",
		mem1 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem10 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem11 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem12 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem13 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem14 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem15 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem16 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem2 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem3 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem4 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem5 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem6 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem7 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem8 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem9 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		OSC_SIM_SETTING => 180000,
		PROGRAM_TIME => 1600000
	  )
	  PORT MAP ( 
		arclk => ufm_arclk,
		ardin => ufm_ardin,
		arshft => ufm_arshft,
		bgpbusy => wire_maxii_ufm_block1_bgpbusy,
		drclk => ufm_drclk,
		drdin => ufm_drdin,
		drdout => wire_maxii_ufm_block1_drdout,
		drshft => ufm_drshft,
		osc => wire_maxii_ufm_block1_osc,
		oscena => ufm_oscena
	  );

 END RTL; --para_altufm_parallel_t9l
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY para IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		nread		: IN STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		nbusy		: OUT STD_LOGIC ;
		osc		: OUT STD_LOGIC 
	);
END para;


ARCHITECTURE RTL OF para IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTUFM_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "access_mode=READ_ONLY;erase_time=500000000;intended_device_family=MAX II;lpm_file=UNUSED;lpm_hint=UNUSED;lpm_type=altufm_parallel;osc_frequency=180000;program_time=1600000;width_address=9;width_data=16;width_ufm_address=9;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC ;



	COMPONENT para_altufm_parallel_t9l
	PORT (
			dataout	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			nread	: IN STD_LOGIC ;
			addr	: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
			data_valid	: OUT STD_LOGIC ;
			nbusy	: OUT STD_LOGIC ;
			osc	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(15 DOWNTO 0);
	data_valid    <= sub_wire1;
	nbusy    <= sub_wire2;
	osc    <= sub_wire3;

	para_altufm_parallel_t9l_component : para_altufm_parallel_t9l
	PORT MAP (
		nread => nread,
		addr => addr,
		dataout => sub_wire0,
		data_valid => sub_wire1,
		nbusy => sub_wire2,
		osc => sub_wire3
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX II"
-- Retrieval info: PRIVATE: OSC_PORT STRING "ON"
-- Retrieval info: CONSTANT: ACCESS_MODE STRING "READ_ONLY"
-- Retrieval info: CONSTANT: ERASE_TIME NUMERIC "500000000"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX II"
-- Retrieval info: CONSTANT: LPM_FILE STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altufm_parallel"
-- Retrieval info: CONSTANT: OSC_FREQUENCY NUMERIC "180000"
-- Retrieval info: CONSTANT: PROGRAM_TIME NUMERIC "1600000"
-- Retrieval info: CONSTANT: WIDTH_ADDRESS NUMERIC "9"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH_UFM_ADDRESS NUMERIC "9"
-- Retrieval info: USED_PORT: addr 0 0 9 0 INPUT NODEFVAL "addr[8..0]"
-- Retrieval info: CONNECT: @addr 0 0 9 0 addr 0 0 9 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: dataout 0 0 16 0 OUTPUT NODEFVAL "dataout[15..0]"
-- Retrieval info: CONNECT: dataout 0 0 16 0 @dataout 0 0 16 0
-- Retrieval info: USED_PORT: nbusy 0 0 0 0 OUTPUT NODEFVAL "nbusy"
-- Retrieval info: CONNECT: nbusy 0 0 0 0 @nbusy 0 0 0 0
-- Retrieval info: USED_PORT: nread 0 0 0 0 INPUT NODEFVAL "nread"
-- Retrieval info: CONNECT: @nread 0 0 0 0 nread 0 0 0 0
-- Retrieval info: USED_PORT: osc 0 0 0 0 OUTPUT NODEFVAL "osc"
-- Retrieval info: CONNECT: osc 0 0 0 0 @osc 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL para.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL para.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL para.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL para_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL para.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL para.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: maxii
